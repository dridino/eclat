-- code generated from the following source code:
--   ../../adrien/stage/vga/test.ecl
--
-- with the following command:
--
--    ./eclat ../../adrien/stage/vga/test.ecl

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.runtime.all;


entity main is
  
  port(signal clk    : in std_logic;
       signal reset  : in std_logic;
       signal run    : in std_logic;
       signal rdy    : out value(0 to 0);
       signal argument : in value(0 to 15);
       signal result : out value(0 to 75));
       
end entity;
architecture rtl of main is

  type t_state is (compute211);
  signal state, \state%next\: t_state;
  type t_state_var229 is (compute222);
  signal state_var229, \state_var229%next\: t_state_var229;
  type t_state_var228 is (compute213, get_pause218, get_wait216, get_wait217, get_wait220);
  signal state_var228, \state_var228%next\: t_state_var228;
  signal \$v227%now\ : value(0 to 0) := (others => '0');
  signal \$v227%next\ : value(0 to 0) := (others => '0');
  signal \$v214%now\ : value(0 to 0) := (others => '0');
  signal \$v214%next\ : value(0 to 0) := (others => '0');
  signal \$496%now\ : value(0 to 21) := (others => '0');
  signal \$496%next\ : value(0 to 21) := (others => '0');
  signal \$499_r_lock%now\ : value(0 to 0) := (others => '0');
  signal \$499_r_lock%next\ : value(0 to 0) := (others => '0');
  signal \rdy221%now\ : value(0 to 0) := (others => '0');
  signal \rdy221%next\ : value(0 to 0) := (others => '0');
  signal \rdy212%now\ : value(0 to 0) := (others => '0');
  signal \rdy212%next\ : value(0 to 0) := (others => '0');
  signal \$482%now\ : value(0 to 14) := (others => '0');
  signal \$482%next\ : value(0 to 14) := (others => '0');
  signal \$490%now\ : value(0 to 14) := (others => '0');
  signal \$490%next\ : value(0 to 14) := (others => '0');
  signal \result209%now\ : value(0 to 75) := (others => '0');
  signal \result209%next\ : value(0 to 75) := (others => '0');
  signal \$v219%now\ : value(0 to 0) := (others => '0');
  signal \$v219%next\ : value(0 to 0) := (others => '0');
  signal \$574%now\ : value(0 to 31) := (others => '0');
  signal \$574%next\ : value(0 to 31) := (others => '0');
  signal \$565%now\ : value(0 to 21) := (others => '0');
  signal \$565%next\ : value(0 to 21) := (others => '0');
  signal \$v215%now\ : value(0 to 0) := (others => '0');
  signal \$v215%next\ : value(0 to 0) := (others => '0');
  signal \rdy210%now\ : value(0 to 0) := (others => '0');
  signal \rdy210%next\ : value(0 to 0) := (others => '0');
  signal \$v207%now\ : value(0 to 43) := (others => '0');
  signal \$v207%next\ : value(0 to 43) := (others => '0');
  signal \$499_r%now\ : value(0 to 31) := (others => '0');
  signal \$499_r%next\ : value(0 to 31) := (others => '0');
  signal \$v225%now\ : value(0 to 0) := (others => '0');
  signal \$v225%next\ : value(0 to 0) := (others => '0');
  signal \$500%now\ : value(0 to 13) := (others => '0');
  signal \$500%next\ : value(0 to 13) := (others => '0');
  signal \$502%now\ : value(0 to 31) := (others => '0');
  signal \$502%next\ : value(0 to 31) := (others => '0');
  signal \$v208%now\ : value(0 to 0) := (others => '0');
  signal \$v208%next\ : value(0 to 0) := (others => '0');
  signal \$v206%now\ : value(0 to 43) := (others => '0');
  signal \$v206%next\ : value(0 to 43) := (others => '0');
  signal \$v224%now\ : value(0 to 0) := (others => '0');
  signal \$v224%next\ : value(0 to 0) := (others => '0');
  
  begin
    process (reset,clk)
        begin
          if reset = '1' then
    \$v227%now\ <= (others => '0');
    \$v214%now\ <= (others => '0');
    \$496%now\ <= (others => '0');
    \$499_r_lock%now\ <= (others => '0');
    \rdy221%now\ <= (others => '0');
    \rdy212%now\ <= (others => '0');
    \$482%now\ <= (others => '0');
    \$490%now\ <= (others => '0');
    \result209%now\ <= (others => '0');
    \$v219%now\ <= (others => '0');
    \$574%now\ <= (others => '0');
    \$565%now\ <= (others => '0');
    \$v215%now\ <= (others => '0');
    \rdy210%now\ <= (others => '0');
    \$v207%now\ <= (others => '0');
    \$499_r%now\ <= (others => '0');
    \$v225%now\ <= (others => '0');
    \$500%now\ <= (others => '0');
    \$502%now\ <= (others => '0');
    \$v208%now\ <= (others => '0');
    \$v206%now\ <= (others => '0');
    \$v224%now\ <= (others => '0');
    state_var229 <= compute222;
    state_var228 <= compute213;
    elsif (rising_edge(clk)) then
    \$v227%now\ <= \$v227%next\;
    \$v214%now\ <= \$v214%next\;
    \$496%now\ <= \$496%next\;
    \$499_r_lock%now\ <= \$499_r_lock%next\;
    \rdy221%now\ <= \rdy221%next\;
    \rdy212%now\ <= \rdy212%next\;
    \$482%now\ <= \$482%next\;
    \$490%now\ <= \$490%next\;
    \result209%now\ <= \result209%next\;
    \$v219%now\ <= \$v219%next\;
    \$574%now\ <= \$574%next\;
    \$565%now\ <= \$565%next\;
    \$v215%now\ <= \$v215%next\;
    \rdy210%now\ <= \rdy210%next\;
    \$v207%now\ <= \$v207%next\;
    \$499_r%now\ <= \$499_r%next\;
    \$v225%now\ <= \$v225%next\;
    \$500%now\ <= \$500%next\;
    \$502%now\ <= \$502%next\;
    \$v208%now\ <= \$v208%next\;
    \$v206%now\ <= \$v206%next\;
    \$v224%now\ <= \$v224%next\;
    state_var229 <= \state_var229%next\;
    state_var228 <= \state_var228%next\;
    state <= \state%next\;
    
    end if;
    end process;
    
    process(argument, clk,state_var229,state_var228, \$v227%now\, \$v214%now\, \$496%now\, \$499_r_lock%now\, \rdy221%now\, \rdy212%now\, \$482%now\, \$490%now\, \result209%now\, \$v219%now\, \$574%now\, \$565%now\, \$v215%now\, \rdy210%now\, \$v207%now\, \$499_r%now\, \$v225%now\, \$500%now\, \$502%now\, \$v208%now\, \$v206%now\, \$v224%now\)
      variable result209 : value(0 to 75) := (others => '0');
      variable \$500\ : value(0 to 13) := (others => '0');
      variable \$v206\, \$v207\ : value(0 to 43) := (others => '0');
      variable \$v224\, \$v208\, \$v225\, rdy210, \$v215\, \$v219\, rdy212, 
               rdy221, \$499_r_lock\, \$v214\, \$v227\ : value(0 to 0) := (others => '0');
      variable \$502\, \$499_r\, \$574\ : value(0 to 31) := (others => '0');
      variable \$490\, \$482\ : value(0 to 14) := (others => '0');
      variable \$565\, \$496\ : value(0 to 21) := (others => '0');
      
    begin
      if run = '1' then
      \$v227\ := \$v227%now\;
      \$v214\ := \$v214%now\;
      \$496\ := \$496%now\;
      \$499_r_lock\ := \$499_r_lock%now\;
      rdy221 := \rdy221%now\;
      rdy212 := \rdy212%now\;
      \$482\ := \$482%now\;
      \$490\ := \$490%now\;
      result209 := \result209%now\;
      \$v219\ := \$v219%now\;
      \$574\ := \$574%now\;
      \$565\ := \$565%now\;
      \$v215\ := \$v215%now\;
      rdy210 := \rdy210%now\;
      \$v207\ := \$v207%now\;
      \$499_r\ := \$499_r%now\;
      \$v225\ := \$v225%now\;
      \$500\ := \$500%now\;
      \$502\ := \$502%now\;
      \$v208\ := \$v208%now\;
      \$v206\ := \$v206%now\;
      \$v224\ := \$v224%now\;
      
      rdy <= "1";
      rdy210 := "0";
      case state is
      when compute211 =>
        rdy210 := eclat_false;
        \$v227\ := eclat_not(rdy212);
        if \$v227\(0) = '1' then
          \$490\ := eclat_true & eclat_true & eclat_true & "0000" & "0000" & "0000";
        end if;
        case state_var228 is
        when get_pause218 =>
          \$499_r_lock\ := eclat_false;
          \$v208\ := eclat_unit;
          if \$499_r_lock\(0) = '1' then
            \state_var228%next\ <= get_wait216;
          else
            \$502\ := \$499_r\;
            eclat_print_int(\$496\(0 to 10));
            
            eclat_print_string(of_string(" "));
            
            eclat_print_int(\$496\(11 to 21));
            
            eclat_print_string(of_string(" "));
            
            \$v215\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false));
            if \$v215\(0) = '1' then
              eclat_print_string(of_string("true"));
              
              \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
              if \$v214\(0) = '1' then
                eclat_print_string(of_string("true"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              else
                eclat_print_string(of_string("false"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              end if;
            else
              eclat_print_string(of_string("false"));
              
              \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
              if \$v214\(0) = '1' then
                eclat_print_string(of_string("true"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              else
                eclat_print_string(of_string("false"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              end if;
            end if;
          end if;
        when get_wait216 =>
          if \$499_r_lock\(0) = '1' then
            \state_var228%next\ <= get_wait216;
          else
            \$502\ := \$499_r\;
            eclat_print_int(\$496\(0 to 10));
            
            eclat_print_string(of_string(" "));
            
            eclat_print_int(\$496\(11 to 21));
            
            eclat_print_string(of_string(" "));
            
            \$v215\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false));
            if \$v215\(0) = '1' then
              eclat_print_string(of_string("true"));
              
              \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
              if \$v214\(0) = '1' then
                eclat_print_string(of_string("true"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              else
                eclat_print_string(of_string("false"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              end if;
            else
              eclat_print_string(of_string("false"));
              
              \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
              if \$v214\(0) = '1' then
                eclat_print_string(of_string("true"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              else
                eclat_print_string(of_string("false"));
                
                eclat_print_newline(eclat_unit);
                
                \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                         eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                \$490\ := eclat_true & \$500\;
                rdy212 := eclat_true;
                \state_var228%next\ <= compute213;
              end if;
            end if;
          end if;
        when get_wait217 =>
          if \$499_r_lock\(0) = '1' then
            \state_var228%next\ <= get_wait217;
          else
            \$499_r_lock\ := eclat_true;
            \$499_r\ := X"0000000" & X"0";
            \state_var228%next\ <= get_pause218;
          end if;
        when get_wait220 =>
          if \$499_r_lock\(0) = '1' then
            \state_var228%next\ <= get_wait220;
          else
            \$574\ := \$499_r\;
            \$v219\ := eclat_if(eclat_eq(\$574\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & 
                       eclat_if(eclat_ge(\$496\(11 to 21) & eclat_vector_get(\$v207\ & X"0000000" & X"1",11)) & 
                       eclat_if(eclat_lt(\$496\(11 to 21) & eclat_add(eclat_vector_get(\$v207\ & X"0000000" & X"1",11) & eclat_vector_get(\$v207\ & X"0000000" & X"3",11))) & 
                       eclat_if(eclat_ge(\$496\(0 to 10) & eclat_vector_get(\$v207\ & X"0000000" & X"0",11)) & eclat_lt(\$496\(0 to 10) & eclat_add(eclat_vector_get(\$v207\ & X"0000000" & X"0",11) & eclat_vector_get(\$v207\ & X"0000000" & X"2",11))) & eclat_false) & eclat_false) & eclat_false) & eclat_false);
            if \$v219\(0) = '1' then
              if \$499_r_lock\(0) = '1' then
                \state_var228%next\ <= get_wait217;
              else
                \$499_r_lock\ := eclat_true;
                \$499_r\ := X"0000000" & X"0";
                \state_var228%next\ <= get_pause218;
              end if;
            else
              \$v208\ := eclat_unit;
              if \$499_r_lock\(0) = '1' then
                \state_var228%next\ <= get_wait216;
              else
                \$502\ := \$499_r\;
                eclat_print_int(\$496\(0 to 10));
                
                eclat_print_string(of_string(" "));
                
                eclat_print_int(\$496\(11 to 21));
                
                eclat_print_string(of_string(" "));
                
                \$v215\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false));
                if \$v215\(0) = '1' then
                  eclat_print_string(of_string("true"));
                  
                  \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
                  if \$v214\(0) = '1' then
                    eclat_print_string(of_string("true"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                    eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                    \$490\ := eclat_true & \$500\;
                    rdy212 := eclat_true;
                    \state_var228%next\ <= compute213;
                  else
                    eclat_print_string(of_string("false"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                    eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                    \$490\ := eclat_true & \$500\;
                    rdy212 := eclat_true;
                    \state_var228%next\ <= compute213;
                  end if;
                else
                  eclat_print_string(of_string("false"));
                  
                  \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
                  if \$v214\(0) = '1' then
                    eclat_print_string(of_string("true"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                    eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                    \$490\ := eclat_true & \$500\;
                    rdy212 := eclat_true;
                    \state_var228%next\ <= compute213;
                  else
                    eclat_print_string(of_string("false"));
                    
                    eclat_print_newline(eclat_unit);
                    
                    \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                    eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                    eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                             eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                    eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                    \$490\ := eclat_true & \$500\;
                    rdy212 := eclat_true;
                    \state_var228%next\ <= compute213;
                  end if;
                end if;
              end if;
            end if;
          end if;
        when compute213 =>
          rdy212 := eclat_false;
          \$v225\ := ""&\$490\(0);
          if \$v225\(0) = '1' then
            \$490\ := eclat_false & \$490\(1 to 14);
            rdy212 := eclat_true;
            \state_var228%next\ <= compute213;
          else
            \$v224\ := eclat_not(rdy221);
            if \$v224\(0) = '1' then
              \$565\ := eclat_sub("00000000000" & "00000000001") & "00000000000";
            end if;
            case state_var229 is
            when compute222 =>
              rdy221 := eclat_false;
              \$565\ := eclat_if(eclat_lt(\$565\(0 to 10) & "01100011111") & eclat_add(\$565\(0 to 10) & "00000000001") & \$565\(11 to 21) & 
                        eclat_if(eclat_lt(\$565\(11 to 21) & "01000001101") & "00000000000" & eclat_add(\$565\(11 to 21) & "00000000001") & "00000000000" & "00000000000"));
              rdy221 := eclat_true;
              \state_var229%next\ <= compute222;
            end case;
            \$565\ := \$565\;
            \$496\ := \$565\;
            \$499_r\ := eclat_sub(X"0000000" & X"0" & X"0000000" & X"1");
            \$v206\ := "00000000000" & "00000000000" & "00000110010" & "00000110010";
            \$v207\ := eclat_vector_get(\$v206\ & X"0000000" & X"0",44);
            if \$499_r_lock\(0) = '1' then
              \state_var228%next\ <= get_wait220;
            else
              \$574\ := \$499_r\;
              \$v219\ := eclat_if(eclat_eq(\$574\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & 
                         eclat_if(eclat_ge(\$496\(11 to 21) & eclat_vector_get(\$v207\ & X"0000000" & X"1",11)) & 
                         eclat_if(eclat_lt(\$496\(11 to 21) & eclat_add(eclat_vector_get(\$v207\ & X"0000000" & X"1",11) & eclat_vector_get(\$v207\ & X"0000000" & X"3",11))) & 
                         eclat_if(eclat_ge(\$496\(0 to 10) & eclat_vector_get(\$v207\ & X"0000000" & X"0",11)) & eclat_lt(\$496\(0 to 10) & eclat_add(eclat_vector_get(\$v207\ & X"0000000" & X"0",11) & eclat_vector_get(\$v207\ & X"0000000" & X"2",11))) & eclat_false) & eclat_false) & eclat_false) & eclat_false);
              if \$v219\(0) = '1' then
                if \$499_r_lock\(0) = '1' then
                  \state_var228%next\ <= get_wait217;
                else
                  \$499_r_lock\ := eclat_true;
                  \$499_r\ := X"0000000" & X"0";
                  \state_var228%next\ <= get_pause218;
                end if;
              else
                \$v208\ := eclat_unit;
                if \$499_r_lock\(0) = '1' then
                  \state_var228%next\ <= get_wait216;
                else
                  \$502\ := \$499_r\;
                  eclat_print_int(\$496\(0 to 10));
                  
                  eclat_print_string(of_string(" "));
                  
                  eclat_print_int(\$496\(11 to 21));
                  
                  eclat_print_string(of_string(" "));
                  
                  \$v215\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false));
                  if \$v215\(0) = '1' then
                    eclat_print_string(of_string("true"));
                    
                    \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
                    if \$v214\(0) = '1' then
                      eclat_print_string(of_string("true"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                      eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                      \$490\ := eclat_true & \$500\;
                      rdy212 := eclat_true;
                      \state_var228%next\ <= compute213;
                    else
                      eclat_print_string(of_string("false"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                      eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                      \$490\ := eclat_true & \$500\;
                      rdy212 := eclat_true;
                      \state_var228%next\ <= compute213;
                    end if;
                  else
                    eclat_print_string(of_string("false"));
                    
                    \$v214\ := eclat_not(eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false));
                    if \$v214\(0) = '1' then
                      eclat_print_string(of_string("true"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                      eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                      \$490\ := eclat_true & \$500\;
                      rdy212 := eclat_true;
                      \state_var228%next\ <= compute213;
                    else
                      eclat_print_string(of_string("false"));
                      
                      eclat_print_newline(eclat_unit);
                      
                      \$500\ := eclat_not(eclat_if(eclat_gt(\$496\(0 to 10) & "00000010000") & eclat_lt(\$496\(0 to 10) & "00001110000") & eclat_false)) & eclat_not(
                      eclat_if(eclat_gt(\$496\(11 to 21) & "00000001010") & eclat_lt(\$496\(11 to 21) & "00000001100") & eclat_false)) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(0 to 3) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(4 to 7) & 
                      eclat_if(eclat_if(eclat_if(eclat_gt(\$496\(0 to 10) & "00000000000") & eclat_lt(\$496\(0 to 10) & "00010100000") & eclat_false) & eclat_true & 
                               eclat_if(eclat_gt(\$496\(11 to 21) & "00000000000") & eclat_lt(\$496\(11 to 21) & "00000101101") & eclat_false)) & "0000" & "0000" & "0000" & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(0 to 3) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(4 to 7) & 
                      eclat_if(eclat_neq(\$502\ & eclat_sub(X"0000000" & X"0" & X"0000000" & X"1")) & "0000" & "0000" & "0000" & "0001" & "0001" & "0001")(8 to 11))(8 to 11);
                      \$490\ := eclat_true & \$500\;
                      rdy212 := eclat_true;
                      \state_var228%next\ <= compute213;
                    end if;
                  end if;
                end if;
              end if;
            end if;
          end if;
        end case;
        \$490\ := \$490\;
        \$482\ := \$490\;
        result209 := argument(0 to 9) & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_true & eclat_false & eclat_false & ""&\$482\(1) & ""&\$482\(2) & \$482\(3 to 6) & \$482\(7 to 10) & \$482\(11 to 14) & eclat_false & eclat_false;
        rdy210 := eclat_true;
        \state%next\ <= compute211;
      end case;\$v227%next\ <= \$v227\;
      \$v214%next\ <= \$v214\;
      \$496%next\ <= \$496\;
      \$499_r_lock%next\ <= \$499_r_lock\;
      \rdy221%next\ <= rdy221;
      \rdy212%next\ <= rdy212;
      \$482%next\ <= \$482\;
      \$490%next\ <= \$490\;
      \result209%next\ <= result209;
      \$v219%next\ <= \$v219\;
      \$574%next\ <= \$574\;
      \$565%next\ <= \$565\;
      \$v215%next\ <= \$v215\;
      \rdy210%next\ <= rdy210;
      \$v207%next\ <= \$v207\;
      \$499_r%next\ <= \$499_r\;
      \$v225%next\ <= \$v225\;
      \$500%next\ <= \$500\;
      \$502%next\ <= \$502\;
      \$v208%next\ <= \$v208\;
      \$v206%next\ <= \$v206\;
      \$v224%next\ <= \$v224\;
      
      
      result <= result209;
      rdy <= rdy210;
      end if;
    end process;
  end architecture;
