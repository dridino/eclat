-- This VHDL was converted from Verilog using the
-- Icarus Verilog VHDL Code Generator 11.0 (stable) ()

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Generated from Verilog module spi_ee_config (spi_ee_config.v:1)
--   ACT_INACT_CTL = 39
--   BW_RATE = 44
--   DATA_FORMAT = 49
--   IDLE = 0
--   IDLE_MSB = 14
--   INI_NUMBER = 11
--   INT_ENABLE = 46
--   INT_MAP = 47
--   INT_SOURCE = 48
--   POWER_CONTROL = 45
--   READ_MODE = 2
--   SI_DataL = 15
--   SO_DataL = 7
--   THRESH_ACT = 36
--   THRESH_FF = 40
--   THRESH_INACT = 37
--   TIME_FF = 41
--   TIME_INACT = 38
--   TRANSFER = 1
--   WRITE_MODE = 0
--   X_HB = 51
--   X_LB = 50
--   Y_HB = 53
--   Y_LB = 52
--   Z_HB = 55
--   Z_LB = 54
entity spi_ee_config is
  port (
    SPI_SDIO : inout std_logic;
    iG_INT2 : in std_logic;
    iRSTN : in std_logic;
    iSPI_CLK : in std_logic;
    iSPI_CLK_OUT : in std_logic;
    data_x : out unsigned(15 downto 0);
    data_y : out unsigned(15 downto 0);
    data_z : out unsigned(15 downto 0);
    oSPI_CLK : out std_logic;
    oSPI_CSN : out std_logic
  );
end entity; 

-- Generated from Verilog module spi_ee_config (spi_ee_config.v:1)
--   ACT_INACT_CTL = 39
--   BW_RATE = 44
--   DATA_FORMAT = 49
--   IDLE = 0
--   IDLE_MSB = 14
--   INI_NUMBER = 11
--   INT_ENABLE = 46
--   INT_MAP = 47
--   INT_SOURCE = 48
--   POWER_CONTROL = 45
--   READ_MODE = 2
--   SI_DataL = 15
--   SO_DataL = 7
--   THRESH_ACT = 36
--   THRESH_FF = 40
--   THRESH_INACT = 37
--   TIME_FF = 41
--   TIME_INACT = 38
--   TRANSFER = 1
--   WRITE_MODE = 0
--   X_HB = 51
--   X_LB = 50
--   Y_HB = 53
--   Y_LB = 52
--   Z_HB = 55
--   Z_LB = 54
architecture from_verilog of spi_ee_config is
  signal clear_status : std_logic;  -- Declared at spi_ee_config.v:42
  signal clear_status_d : unsigned(3 downto 0);  -- Declared at spi_ee_config.v:43
  signal high_byte : std_logic;  -- Declared at spi_ee_config.v:40
  signal high_byte_d : std_logic;  -- Declared at spi_ee_config.v:44
  signal ini_index : unsigned(3 downto 0);  -- Declared at spi_ee_config.v:32
  signal low_byte_data : unsigned(7 downto 0);  -- Declared at spi_ee_config.v:38
  signal p2s_data : unsigned(15 downto 0);  -- Declared at spi_ee_config.v:34
  signal read_back : std_logic;  -- Declared at spi_ee_config.v:41
  signal read_back_d : std_logic;  -- Declared at spi_ee_config.v:44
  signal read_idle_count : unsigned(14 downto 0);  -- Declared at spi_ee_config.v:45
  signal read_ready : std_logic;  -- Declared at spi_ee_config.v:42
  signal s2p_data : unsigned(7 downto 0);  -- Declared at spi_ee_config.v:37
  signal spi_end : std_logic;  -- Declared at spi_ee_config.v:36
  signal spi_go : std_logic;  -- Declared at spi_ee_config.v:35
  signal spi_state : std_logic;  -- Declared at spi_ee_config.v:39
  signal write_data : unsigned(13 downto 0);  -- Declared at spi_ee_config.v:33
  -- ajout
  signal read_idx : integer range 0 to 2; -- 0 -> x; 1 -> y; 2 -> z

  component spi_controller is
    port (
      SPI_SDIO : inout std_logic;
      iP2S_DATA : in unsigned(15 downto 0);
      iRSTN : in std_logic;
      iSPI_CLK : in std_logic;
      iSPI_CLK_OUT : in std_logic;
      iSPI_GO : in std_logic;
      oS2P_DATA : out unsigned(7 downto 0);
      oSPI_CLK : out std_logic;
      oSPI_CSN : out std_logic;
      oSPI_END : buffer std_logic
    );
  end component;
  signal oSPI_CLK_Readable : std_logic;  -- Needed to connect outputs
  signal oSPI_CSN_Readable : std_logic;  -- Needed to connect outputs
begin
  oSPI_CLK <= oSPI_CLK_Readable;
  oSPI_CSN <= oSPI_CSN_Readable;
  
  -- Generated from instantiation at spi_ee_config.v:50
  u_spi_controller: spi_controller
    port map (
      SPI_SDIO => SPI_SDIO,
      iP2S_DATA => p2s_data,
      iRSTN => iRSTN,
      iSPI_CLK => iSPI_CLK,
      iSPI_CLK_OUT => iSPI_CLK_OUT,
      iSPI_GO => spi_go,
      oS2P_DATA => s2p_data,
      oSPI_CLK => oSPI_CLK_Readable,
      oSPI_CSN => oSPI_CSN_Readable,
      oSPI_END => spi_end
    );
  
  -- Generated from always process in spi_ee_config (spi_ee_config.v:66)
  process (ini_index) is
  begin
    case ini_index is
      when X"0" =>
        write_data <= "10010000100000";
      when X"1" =>
        write_data <= "10010100000011";
      when X"2" =>
        write_data <= "10011000000001";
      when X"3" =>
        write_data <= "10011101111111";
      when X"4" =>
        write_data <= "10100000001001";
      when X"5" =>
        write_data <= "10100101000110";
      when X"6" =>
        write_data <= "10110000001001";
      when X"7" =>
        write_data <= "10111000010000";
      when X"8" =>
        write_data <= "10111100010000";
      when X"9" =>
        write_data <= "11000101000000";
      when others =>
        write_data <= "10110100001000";
    end case;
  end process;
  
  -- Generated from always process in spi_ee_config (spi_ee_config.v:81)
  process (iRSTN, iSPI_CLK) is
  begin
    if (not iRSTN) = '1' then
      ini_index <= X"0";
      spi_go <= '0';
      spi_state <= '0';
      read_idle_count <= "000000000000000";
      high_byte <= '0';
      read_idx <= 1;
      read_back <= '0';
      clear_status <= '0';
    elsif rising_edge(iSPI_CLK) then
      if ini_index < X"b" then
        case spi_state is
          when '0' =>
            p2s_data <= "00" & write_data;
            spi_go <= '1';
            spi_state <= '1';
          when '1' =>
            if spi_end = '1' then
              ini_index <= ini_index + X"1";
              spi_go <= '0';
              spi_state <= '0';
            end if;
          when others =>
            null;
        end case;
      else
        case spi_state is
          when '0' =>
            read_idle_count <= read_idle_count + "000000000000001";
            if high_byte = '1' then
              case read_idx is
                when 0 => p2s_data(8 + 7 downto 8) <= "10110011"; -- READMODE(2) & X_HB(6)
                when 1 => p2s_data(8 + 7 downto 8) <= "10110101"; -- READMODE(2) & Y_HB(6)
                when 2 => p2s_data(8 + 7 downto 8) <= "10110111"; -- READMODE(2) & Z_HB(6)
                when others => null;
              end case;
              read_back <= '1';
            else
              if read_ready = '1' then
                case read_idx is
                  when 0 => p2s_data(8 + 7 downto 8) <= "10110010"; -- READMODE(2) & X_LB(6)
                  when 1 => p2s_data(8 + 7 downto 8) <= "10110100"; -- READMODE(2) & Y_LB(6)
                  when 2 => p2s_data(8 + 7 downto 8) <= "10110110"; -- READMODE(2) & Z_LB(6)
                  when others => null;
                end case;
                read_back <= '1';
              else
                if (((not clear_status_d(3)) = '1') and (iG_INT2 = '1')) or (read_idle_count(14) = '1') then
                  p2s_data(8 + 7 downto 8) <= X"b0";
                  clear_status <= '1';
                end if;
              end if;
            end if;
            if (((high_byte = '1') or (read_ready = '1')) or (read_idle_count(14) = '1')) or (((not clear_status_d(3)) = '1') and (iG_INT2 = '1')) then
              spi_go <= '1';
              spi_state <= '1';
            end if;
            if read_back_d = '1' then
              if high_byte_d = '1' then
                case read_idx is
                  when 0 => data_z <= s2p_data & low_byte_data;
                  when 1 => data_x <= s2p_data & low_byte_data;
                  when 2 => data_y <= s2p_data & low_byte_data;
                  when others => null;
                end case;
              else
                low_byte_data <= s2p_data;
              end if;
            end if;
          when '1' =>
            if spi_end = '1' then
              spi_go <= '0';
              spi_state <= '0';
              if read_back = '1' then
                read_back <= '0';
                if high_byte = '1' then
                  if read_idx = 2 then
                    read_idx <= 0;
                  else
                    read_idx <= read_idx + 1;
                  end if;
                end if;
                high_byte <= not high_byte;
                read_ready <= '0';
              else
                clear_status <= '0';
                read_ready <= s2p_data(6);
                read_idle_count <= "000000000000000";
              end if;
            end if;
          when others =>
            null;
        end case;
      end if;
    end if;
  end process;
  
  -- Generated from always process in spi_ee_config (spi_ee_config.v:170)
  process (iRSTN, iSPI_CLK) is
  begin
    if (not iRSTN) = '1' then
      high_byte_d <= '0';
      read_back_d <= '0';
      clear_status_d <= X"0";
    elsif rising_edge(iSPI_CLK) then
      high_byte_d <= high_byte;
      read_back_d <= read_back;
      clear_status_d <= clear_status_d(0 + 2 downto 0) & clear_status;
    end if;
  end process;
end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Generated from Verilog module spi_controller (spi_controller.v:1)
--   ACT_INACT_CTL = 39
--   BW_RATE = 44
--   DATA_FORMAT = 49
--   IDLE = 0
--   IDLE_MSB = 14
--   INI_NUMBER = 11
--   INT_ENABLE = 46
--   INT_MAP = 47
--   INT_SOURCE = 48
--   POWER_CONTROL = 45
--   READ_MODE = 2
--   SI_DataL = 15
--   SO_DataL = 7
--   THRESH_ACT = 36
--   THRESH_FF = 40
--   THRESH_INACT = 37
--   TIME_FF = 41
--   TIME_INACT = 38
--   TRANSFER = 1
--   WRITE_MODE = 0
--   X_HB = 51
--   X_LB = 50
--   Y_HB = 53
--   Y_LB = 52
--   Z_HB = 55
--   Z_LB = 54
entity spi_controller is
  port (
    SPI_SDIO : inout std_logic;
    iP2S_DATA : in unsigned(15 downto 0);
    iRSTN : in std_logic;
    iSPI_CLK : in std_logic;
    iSPI_CLK_OUT : in std_logic;
    iSPI_GO : in std_logic;
    oS2P_DATA : out unsigned(7 downto 0);
    oSPI_CLK : out std_logic;
    oSPI_CSN : out std_logic;
    oSPI_END : buffer std_logic
  );
end entity; 

-- Generated from Verilog module spi_controller (spi_controller.v:1)
--   ACT_INACT_CTL = 39
--   BW_RATE = 44
--   DATA_FORMAT = 49
--   IDLE = 0
--   IDLE_MSB = 14
--   INI_NUMBER = 11
--   INT_ENABLE = 46
--   INT_MAP = 47
--   INT_SOURCE = 48
--   POWER_CONTROL = 45
--   READ_MODE = 2
--   SI_DataL = 15
--   SO_DataL = 7
--   THRESH_ACT = 36
--   THRESH_FF = 40
--   THRESH_INACT = 37
--   TIME_FF = 41
--   TIME_INACT = 38
--   TRANSFER = 1
--   WRITE_MODE = 0
--   X_HB = 51
--   X_LB = 50
--   Y_HB = 53
--   Y_LB = 52
--   Z_HB = 55
--   Z_LB = 54
architecture from_verilog of spi_controller is
  signal oS2P_DATA_Reg : unsigned(7 downto 0);
  signal tmp_ivl_13 : std_logic;  -- Temporary created at spi_controller.v:46
  signal tmp_ivl_15 : std_logic;  -- Temporary created at spi_controller.v:46
  signal tmp_ivl_17 : std_logic;  -- Temporary created at spi_controller.v:46
  signal tmp_ivl_19 : std_logic;  -- Temporary created at spi_controller.v:46
  signal read_mode : std_logic;  -- Declared at spi_controller.v:34
  signal spi_count : unsigned(3 downto 0);  -- Declared at spi_controller.v:36
  signal spi_count_en : std_logic;  -- Declared at spi_controller.v:35
  signal write_address : std_logic;  -- Declared at spi_controller.v:34
  
  function Reduce_OR(X : std_logic_vector) return std_logic is
    variable R : std_logic := '0';
  begin
    for I in X'Range loop
      R := X(I) or R;
    end loop;
    return R;
  end function;
begin
  oS2P_DATA <= oS2P_DATA_Reg;
  oSPI_CSN <= not iSPI_GO;
  tmp_ivl_15 <= tmp_ivl_13 or write_address;
  tmp_ivl_17 <= spi_count_en and tmp_ivl_15;
  read_mode <= iP2S_DATA(15);
  write_address <= spi_count(3);
  oSPI_END <= not Reduce_OR(std_logic_vector(spi_count));
  oSPI_CLK <= iSPI_CLK_OUT when spi_count_en = '1' else '1';
  tmp_ivl_13 <= not read_mode;
  tmp_ivl_19 <= iP2S_DATA(To_Integer(spi_count));
  SPI_SDIO <= tmp_ivl_19 when tmp_ivl_17 = '1' else 'Z';
  
  -- Generated from always process in spi_controller (spi_controller.v:48)
  process (iRSTN, iSPI_CLK) is
  begin
    if (not iRSTN) = '1' then
      spi_count_en <= '0';
      spi_count <= X"f";
    elsif rising_edge(iSPI_CLK) then
      if oSPI_END = '1' then
        spi_count_en <= '0';
      else
        if iSPI_GO = '1' then
          spi_count_en <= '1';
        end if;
      end if;
      if (not spi_count_en) = '1' then
        spi_count <= X"f";
      else
        spi_count <= spi_count - X"1";
      end if;
      if (read_mode = '1') and ((not write_address) = '1') then
        oS2P_DATA_Reg <= oS2P_DATA_Reg(0 + 6 downto 0) & SPI_SDIO;
      end if;
    end if;
  end process;
end architecture;

